`ifndef SSEMI_TIMESCALE_VH
`define SSEMI_TIMESCALE_VH

//=============================================================================
// Common Timescale Definition
//=============================================================================
// Description: Standard timescale for SSEMI ADC Decimator IP
// Author:      SSEMI Development Team
// Date:        2025-08-30T18:32:01Z
// License:     Apache-2.0
//=============================================================================

`timescale 1ns/1ps

`endif // SSEMI_TIMESCALE_VH
